��/ /   ! !   D o   n o t   e d i t   -   a u t o - g e n e r a t e d   ! !  
  
 / * - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
     m o d u l e n a m e   :   a p b _ p l i c _ r e g s  
     g e n e r a t e d   b y   A n t o n   D u m a s   o n   1 7 / 0 1 / 2 0 2 2   0 0 : 5 5 : 2 4   w i t h   0 . 1   A l p h a  
  
     d e s c r i p t i o n :   P L I C   A d d r e s s   M a p  
 - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - * /  
  
 m o d u l e   a p b _ p l i c _ r e g s  
 (  
     / /   p o r t   p r i o   ( A c c e s s . R W )  
     i n p u t     l o g i c   [ 7 0 : 0 ] [ 2 : 0 ]   p r i o _ i ,  
     o u t p u t   l o g i c   [ 7 0 : 0 ]   p r i o _ r e _ o ,  
     o u t p u t   l o g i c   [ 7 0 : 0 ] [ 2 : 0 ]   p r i o _ o ,  
     o u t p u t   l o g i c   [ 7 0 : 0 ]   p r i o _ w e _ o ,  
  
     / /   p o r t   i p   ( A c c e s s . R O )  
     i n p u t     l o g i c   [ 7 0 : 0 ]   i p _ i ,  
     o u t p u t   l o g i c     i p _ r e _ o ,  
  
     / /   p o r t   i e   ( A c c e s s . R W )  
     i n p u t     l o g i c   [ 1 : 0 ] [ 7 0 : 0 ]   i e _ i ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   i e _ r e _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ] [ 7 0 : 0 ]   i e _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   i e _ w e _ o ,  
  
     / /   p o r t   t h r e s h o l d   ( A c c e s s . R W )  
     i n p u t     l o g i c   [ 1 : 0 ] [ 2 : 0 ]   t h r e s h o l d _ i ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   t h r e s h o l d _ r e _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ] [ 2 : 0 ]   t h r e s h o l d _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   t h r e s h o l d _ w e _ o ,  
  
     / /   p o r t   c c   ( A c c e s s . R W )  
     i n p u t     l o g i c   [ 1 : 0 ] [ 6 : 0 ]   c c _ i ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   c c _ r e _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ] [ 6 : 0 ]   c c _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   c c _ w e _ o ,  
  
  
     / /   A P B 3   i n t e r f a c e  
     i n p u t     l o g i c   [ 3 1 : 0 ]   p a d d r _ i ,  
     i n p u t     l o g i c                 p s e l _ i ,  
     i n p u t     l o g i c                 p e n a b l e _ i ,  
     i n p u t     l o g i c                 p w r i t e _ i ,  
     i n p u t     l o g i c   [ 3 1 : 0 ]   p w d a t a _ i ,  
     o u t p u t   l o g i c   [ 3 1 : 0 ]   p r d a t a _ o ,  
     o u t p u t   l o g i c                 p r e a d y _ o ,  
     o u t p u t   l o g i c                 p s l v e r r _ o  
 ) ;  
  
     / /   c o m b i n a t o r i a l   r e g i s t e r   m u x  
     a l w a y s _ c o m b   b e g i n   :   b e g i n _ g e n _ r e g _ m u x _ a p b _ p l i c _ r e g s  
         / /   a p b 3   b u s   d e f a u l t s  
         p r e a d y _ o     =   1 ' b 1 ;   / /   s l a v e   i s   a l w a y s   r e a d y  
         p r d a t a _ o     =       ' 0 ;  
         p s l v e r r _ o   =       ' 0 ;  
         / /   r e g   p o r t s   d e f a u l t s  
         / /   r e g   p r i o   d e f a u l t s  
         p r i o _ o         =   ' 0 ;  
         p r i o _ w e _ o   =   ' 0 ;  
         p r i o _ r e _ o   =   ' 0 ;  
         / /   r e g   i p   d e f a u l t s  
         i p _ r e _ o   =   ' 0 ;  
         / /   r e g   i e   d e f a u l t s  
         i e _ o         =   ' 0 ;  
         i e _ w e _ o   =   ' 0 ;  
         i e _ r e _ o   =   ' 0 ;  
         / /   r e g   t h r e s h o l d   d e f a u l t s  
         t h r e s h o l d _ o         =   ' 0 ;  
         t h r e s h o l d _ w e _ o   =   ' 0 ;  
         t h r e s h o l d _ r e _ o   =   ' 0 ;  
         / /   r e g   c c   d e f a u l t s  
         c c _ o         =   ' 0 ;  
         c c _ w e _ o   =   ' 0 ;  
         c c _ r e _ o   =   ' 0 ;  
         / /   a p b 3   b u s   w r i t e   l o g i c  
         i f   ( p s e l _ i   &   p e n a b l e _ i )   b e g i n  
             i f   ( p w r i t e _ i )   b e g i n  
                 u n i q u e   c a s e ( p a d d r _ i )  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 0   :   b e g i n  
                         p r i o _ i [ 0 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 4   :   b e g i n  
                         p r i o _ i [ 1 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 8   :   b e g i n  
                         p r i o _ i [ 2 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 c   :   b e g i n  
                         p r i o _ i [ 3 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 0   :   b e g i n  
                         p r i o _ i [ 4 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 4   :   b e g i n  
                         p r i o _ i [ 5 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 8   :   b e g i n  
                         p r i o _ i [ 6 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 c   :   b e g i n  
                         p r i o _ i [ 7 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 0   :   b e g i n  
                         p r i o _ i [ 8 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 4   :   b e g i n  
                         p r i o _ i [ 9 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 8   :   b e g i n  
                         p r i o _ i [ 1 0 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 c   :   b e g i n  
                         p r i o _ i [ 1 1 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 0   :   b e g i n  
                         p r i o _ i [ 1 2 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 4   :   b e g i n  
                         p r i o _ i [ 1 3 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 8   :   b e g i n  
                         p r i o _ i [ 1 4 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 c   :   b e g i n  
                         p r i o _ i [ 1 5 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 0   :   b e g i n  
                         p r i o _ i [ 1 6 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 4   :   b e g i n  
                         p r i o _ i [ 1 7 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 8   :   b e g i n  
                         p r i o _ i [ 1 8 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 c   :   b e g i n  
                         p r i o _ i [ 1 9 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 0   :   b e g i n  
                         p r i o _ i [ 2 0 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 4   :   b e g i n  
                         p r i o _ i [ 2 1 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 8   :   b e g i n  
                         p r i o _ i [ 2 2 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 c   :   b e g i n  
                         p r i o _ i [ 2 3 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 0   :   b e g i n  
                         p r i o _ i [ 2 4 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 4   :   b e g i n  
                         p r i o _ i [ 2 5 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 8   :   b e g i n  
                         p r i o _ i [ 2 6 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 c   :   b e g i n  
                         p r i o _ i [ 2 7 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 0   :   b e g i n  
                         p r i o _ i [ 2 8 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 4   :   b e g i n  
                         p r i o _ i [ 2 9 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 8   :   b e g i n  
                         p r i o _ i [ 3 0 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 c   :   b e g i n  
                         p r i o _ i [ 3 1 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 8 0   :   b e g i n  
                         p r i o _ i [ 3 2 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 8 4   :   b e g i n  
                         p r i o _ i [ 3 3 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 8 8   :   b e g i n  
                         p r i o _ i [ 3 4 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 8 c   :   b e g i n  
                         p r i o _ i [ 3 5 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 9 0   :   b e g i n  
                         p r i o _ i [ 3 6 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 9 4   :   b e g i n  
                         p r i o _ i [ 3 7 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 9 8   :   b e g i n  
                         p r i o _ i [ 3 8 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 9 c   :   b e g i n  
                         p r i o _ i [ 3 9 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 a 0   :   b e g i n  
                         p r i o _ i [ 4 0 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 a 4   :   b e g i n  
                         p r i o _ i [ 4 1 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 a 8   :   b e g i n  
                         p r i o _ i [ 4 2 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 a c   :   b e g i n  
                         p r i o _ i [ 4 3 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 b 0   :   b e g i n  
                         p r i o _ i [ 4 4 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 b 4   :   b e g i n  
                         p r i o _ i [ 4 5 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 b 8   :   b e g i n  
                         p r i o _ i [ 4 6 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 b c   :   b e g i n  
                         p r i o _ i [ 4 7 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 c 0   :   b e g i n  
                         p r i o _ i [ 4 8 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 c 4   :   b e g i n  
                         p r i o _ i [ 4 9 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 c 8   :   b e g i n  
                         p r i o _ i [ 5 0 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 c c   :   b e g i n  
                         p r i o _ i [ 5 1 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 d 0   :   b e g i n  
                         p r i o _ i [ 5 2 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 d 4   :   b e g i n  
                         p r i o _ i [ 5 3 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 d 8   :   b e g i n  
                         p r i o _ i [ 5 4 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 d c   :   b e g i n  
                         p r i o _ i [ 5 5 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 e 0   :   b e g i n  
                         p r i o _ i [ 5 6 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 e 4   :   b e g i n  
                         p r i o _ i [ 5 7 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 e 8   :   b e g i n  
                         p r i o _ i [ 5 8 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 e c   :   b e g i n  
                         p r i o _ i [ 5 9 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 f 0   :   b e g i n  
                         p r i o _ i [ 6 0 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 f 4   :   b e g i n  
                         p r i o _ i [ 6 1 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 f 8   :   b e g i n  
                         p r i o _ i [ 6 2 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 f c   :   b e g i n  
                         p r i o _ i [ 6 3 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 0 0   :   b e g i n  
                         p r i o _ i [ 6 4 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 0 4   :   b e g i n  
                         p r i o _ i [ 6 5 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 0 8   :   b e g i n  
                         p r i o _ i [ 6 6 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 0 c   :   b e g i n  
                         p r i o _ i [ 6 7 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 1 0   :   b e g i n  
                         p r i o _ i [ 6 8 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 1 4   :   b e g i n  
                         p r i o _ i [ 6 9 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 1 8   :   b e g i n  
                         p r i o _ i [ 7 0 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 7 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 0 0   :   b e g i n  
                         i e _ i [ 0 ] [ 3 1 : 0 ]   =   p w d a t a _ i [ 3 1 : 0 ] ;  
                         i e _ w e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 8 0   :   b e g i n  
                         i e _ i [ 1 ] [ 3 1 : 0 ]   =   p w d a t a _ i [ 3 1 : 0 ] ;  
                         i e _ w e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 0 4   :   b e g i n  
                         i e _ i [ 0 ] [ 6 3 : 3 2 ]   =   p w d a t a _ i [ 3 1 : 0 ] ;  
                         i e _ w e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 8 4   :   b e g i n  
                         i e _ i [ 1 ] [ 6 3 : 3 2 ]   =   p w d a t a _ i [ 3 1 : 0 ] ;  
                         i e _ w e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 0 8   :   b e g i n  
                         i e _ i [ 0 ] [ 7 0 : 6 4 ]   =   p w d a t a _ i [ 6 : 0 ] ;  
                         i e _ w e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 8 8   :   b e g i n  
                         i e _ i [ 1 ] [ 7 0 : 6 4 ]   =   p w d a t a _ i [ 6 : 0 ] ;  
                         i e _ w e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   t h r e s h o l d  
                     3 2 ' h c 2 0 0 0 0 0   :   b e g i n  
                         t h r e s h o l d _ i [ 0 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         t h r e s h o l d _ w e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   t h r e s h o l d  
                     3 2 ' h c 2 0 1 0 0 0   :   b e g i n  
                         t h r e s h o l d _ i [ 1 ] [ 2 : 0 ]   =   p w d a t a _ i [ 2 : 0 ] ;  
                         t h r e s h o l d _ w e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   c c  
                     3 2 ' h c 2 0 0 0 0 4   :   b e g i n  
                         c c _ i [ 0 ] [ 6 : 0 ]   =   p w d a t a _ i [ 6 : 0 ] ;  
                         c c _ w e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   c c  
                     3 2 ' h c 2 0 0 0 0 8   :   b e g i n  
                         c c _ i [ 1 ] [ 6 : 0 ]   =   p w d a t a _ i [ 6 : 0 ] ;  
                         c c _ w e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     d e f a u l t :   b e g i n    
                         p s l v e r r _ o   =   1 ' b 1 ;  
                     e n d  
                 e n d c a s e  
             e n d   e l s e   b e g i n  
                 u n i q u e   c a s e ( p a d d r _ i )  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 1 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 2 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 3 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 4 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 5 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 6 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 7 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 8 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 9 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 1 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 1 1 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 1 2 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 1 3 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 1 4 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 1 5 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 1 6 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 1 7 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 1 8 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 1 9 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 2 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 2 1 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 2 2 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 2 3 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 2 4 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 2 5 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 2 6 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 2 7 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 2 8 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 2 9 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 3 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 3 1 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 8 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 3 2 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 8 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 3 3 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 8 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 3 4 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 8 c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 3 5 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 9 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 3 6 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 9 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 3 7 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 9 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 3 8 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 9 c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 3 9 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 a 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 4 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 a 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 4 1 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 a 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 4 2 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 a c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 4 3 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 b 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 4 4 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 b 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 4 5 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 b 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 4 6 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 b c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 4 7 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 c 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 4 8 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 c 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 4 9 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 c 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 5 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 c c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 5 1 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 d 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 5 2 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 d 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 5 3 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 d 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 5 4 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 d c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 5 5 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 e 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 5 6 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 e 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 5 7 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 e 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 5 8 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 e c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 5 9 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 f 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 6 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 f 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 6 1 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 f 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 6 2 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 f c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 6 3 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 0 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 6 4 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 0 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 6 5 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 0 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 6 6 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 0 c   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 6 7 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 1 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 6 8 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 1 4   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 6 9 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 1 1 8   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   p r i o _ o [ 7 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 7 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i p  
                     3 2 ' h c 0 0 1 0 0 0   :   b e g i n  
                         p r d a t a _ o [ 3 1 : 0 ]   =   i p _ o [ 3 1 : 0 ] ;  
                         i p _ r e _ o   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i p  
                     3 2 ' h c 0 0 1 0 0 4   :   b e g i n  
                         p r d a t a _ o [ 3 1 : 0 ]   =   i p _ o [ 6 3 : 3 2 ] ;  
                         i p _ r e _ o   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i p  
                     3 2 ' h c 0 0 1 0 0 8   :   b e g i n  
                         p r d a t a _ o [ 6 : 0 ]   =   i p _ o [ 7 0 : 6 4 ] ;  
                         i p _ r e _ o   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 0 0   :   b e g i n  
                         p r d a t a _ o [ 3 1 : 0 ]   =   i e _ o [ 0 ] [ 3 1 : 0 ] ;  
                         i e _ r e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 8 0   :   b e g i n  
                         p r d a t a _ o [ 3 1 : 0 ]   =   i e _ o [ 1 ] [ 3 1 : 0 ] ;  
                         i e _ r e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 0 4   :   b e g i n  
                         p r d a t a _ o [ 3 1 : 0 ]   =   i e _ o [ 0 ] [ 6 3 : 3 2 ] ;  
                         i e _ r e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 8 4   :   b e g i n  
                         p r d a t a _ o [ 3 1 : 0 ]   =   i e _ o [ 1 ] [ 6 3 : 3 2 ] ;  
                         i e _ r e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 0 8   :   b e g i n  
                         p r d a t a _ o [ 6 : 0 ]   =   i e _ o [ 0 ] [ 7 0 : 6 4 ] ;  
                         i e _ r e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 8 8   :   b e g i n  
                         p r d a t a _ o [ 6 : 0 ]   =   i e _ o [ 1 ] [ 7 0 : 6 4 ] ;  
                         i e _ r e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   t h r e s h o l d  
                     3 2 ' h c 2 0 0 0 0 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   t h r e s h o l d _ o [ 0 ] [ 2 : 0 ] ;  
                         t h r e s h o l d _ r e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   t h r e s h o l d  
                     3 2 ' h c 2 0 1 0 0 0   :   b e g i n  
                         p r d a t a _ o [ 2 : 0 ]   =   t h r e s h o l d _ o [ 1 ] [ 2 : 0 ] ;  
                         t h r e s h o l d _ r e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   c c  
                     3 2 ' h c 2 0 0 0 0 4   :   b e g i n  
                         p r d a t a _ o [ 6 : 0 ]   =   c c _ o [ 0 ] [ 6 : 0 ] ;  
                         c c _ r e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   c c  
                     3 2 ' h c 2 0 0 0 0 8   :   b e g i n  
                         p r d a t a _ o [ 6 : 0 ]   =   c c _ o [ 1 ] [ 6 : 0 ] ;  
                         c c _ r e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     d e f a u l t :   b e g i n    
                         p s l v e r r _ o   =   1 ' b 1 ;  
                     e n d  
                 e n d c a s e  
             e n d  
         e n d  
     e n d   :   e n d _ g e n _ r e g _ m u x _ a p b _ p l i c _ r e g s  
 e n d m o d u l e  
  
 