��/ /   ! !   D o   n o t   e d i t   -   a u t o - g e n e r a t e d   ! !  
  
 / * - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
     m o d u l e n a m e   :   p l i c _ r e g s  
     g e n e r a t e d   b y   A n t o n   D u m a s   o n   1 7 / 0 1 / 2 0 2 2   0 9 : 3 4 : 0 1   w i t h   0 . 1   A l p h a  
  
     d e s c r i p t i o n :   P L I C   A d d r e s s   M a p  
 - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - * /  
  
 m o d u l e   p l i c _ r e g s  
 (  
     / /   p o r t   p r i o   ( A c c e s s . R W )  
     i n p u t     l o g i c   [ 3 0 : 0 ] [ 2 : 0 ]   p r i o _ i ,  
     o u t p u t   l o g i c   [ 3 0 : 0 ]   p r i o _ r e _ o ,  
     o u t p u t   l o g i c   [ 3 0 : 0 ] [ 2 : 0 ]   p r i o _ o ,  
     o u t p u t   l o g i c   [ 3 0 : 0 ]   p r i o _ w e _ o ,  
  
     / /   p o r t   i p   ( A c c e s s . R O )  
     i n p u t     l o g i c   [ 3 0 : 0 ]   i p _ i ,  
     o u t p u t   l o g i c     i p _ r e _ o ,  
  
     / /   p o r t   i e   ( A c c e s s . R W )  
     i n p u t     l o g i c   [ 1 : 0 ] [ 3 0 : 0 ]   i e _ i ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   i e _ r e _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ] [ 3 0 : 0 ]   i e _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   i e _ w e _ o ,  
  
     / /   p o r t   t h r e s h o l d   ( A c c e s s . R W )  
     i n p u t     l o g i c   [ 1 : 0 ] [ 2 : 0 ]   t h r e s h o l d _ i ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   t h r e s h o l d _ r e _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ] [ 2 : 0 ]   t h r e s h o l d _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   t h r e s h o l d _ w e _ o ,  
  
     / /   p o r t   c c   ( A c c e s s . R W )  
     i n p u t     l o g i c   [ 1 : 0 ] [ 4 : 0 ]   c c _ i ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   c c _ r e _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ] [ 4 : 0 ]   c c _ o ,  
     o u t p u t   l o g i c   [ 1 : 0 ]   c c _ w e _ o ,  
  
  
     / /   B u s   I n t e r f a c e  
     i n p u t     r e g _ i n t f : : r e g _ i n t f _ r e q _ a 3 2 _ d 3 2   r e q _ i ,  
     o u t p u t   r e g _ i n t f : : r e g _ i n t f _ r e s p _ d 3 2         r e s p _ o  
 ) ;  
  
     / /   c o m b i n a t o r i a l   r e g i s t e r   m u x  
     a l w a y s _ c o m b   b e g i n   :   b e g i n _ g e n _ r e g _ m u x _ p l i c _ r e g s  
         / /   r e g   b u s   d e f a u l t s  
         r e s p _ o . r e a d y   =   1 ' b 1 ;   / /   s l a v e   i s   a l w a y s   r e a d y  
         r e s p _ o . r d a t a   =       ' 0 ;  
         r e s p _ o . e r r o r   =       ' 0 ;  
         / /   r e g   p o r t s   d e f a u l t s  
         / /   r e g   p r i o   d e f a u l t s  
         p r i o _ o         =   ' 0 ;  
         p r i o _ w e _ o   =   ' 0 ;  
         p r i o _ r e _ o   =   ' 0 ;  
         / /   r e g   i p   d e f a u l t s  
         i p _ r e _ o   =   ' 0 ;  
         / /   r e g   i e   d e f a u l t s  
         i e _ o         =   ' 0 ;  
         i e _ w e _ o   =   ' 0 ;  
         i e _ r e _ o   =   ' 0 ;  
         / /   r e g   t h r e s h o l d   d e f a u l t s  
         t h r e s h o l d _ o         =   ' 0 ;  
         t h r e s h o l d _ w e _ o   =   ' 0 ;  
         t h r e s h o l d _ r e _ o   =   ' 0 ;  
         / /   r e g   c c   d e f a u l t s  
         c c _ o         =   ' 0 ;  
         c c _ w e _ o   =   ' 0 ;  
         c c _ r e _ o   =   ' 0 ;  
         / /   r e g   b u s   w r i t e   l o g i c  
         i f   ( r e q _ i . v a l i d )   b e g i n  
             i f   ( r e q _ i . w r i t e )   b e g i n  
                 u n i q u e   c a s e ( r e q _ i . a d d r )  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 0   :   b e g i n  
                         p r i o _ i [ 0 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 4   :   b e g i n  
                         p r i o _ i [ 1 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 8   :   b e g i n  
                         p r i o _ i [ 2 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 c   :   b e g i n  
                         p r i o _ i [ 3 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 0   :   b e g i n  
                         p r i o _ i [ 4 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 4   :   b e g i n  
                         p r i o _ i [ 5 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 8   :   b e g i n  
                         p r i o _ i [ 6 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 c   :   b e g i n  
                         p r i o _ i [ 7 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 0   :   b e g i n  
                         p r i o _ i [ 8 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 4   :   b e g i n  
                         p r i o _ i [ 9 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 8   :   b e g i n  
                         p r i o _ i [ 1 0 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 c   :   b e g i n  
                         p r i o _ i [ 1 1 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 0   :   b e g i n  
                         p r i o _ i [ 1 2 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 4   :   b e g i n  
                         p r i o _ i [ 1 3 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 8   :   b e g i n  
                         p r i o _ i [ 1 4 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 c   :   b e g i n  
                         p r i o _ i [ 1 5 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 0   :   b e g i n  
                         p r i o _ i [ 1 6 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 4   :   b e g i n  
                         p r i o _ i [ 1 7 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 8   :   b e g i n  
                         p r i o _ i [ 1 8 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 c   :   b e g i n  
                         p r i o _ i [ 1 9 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 1 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 0   :   b e g i n  
                         p r i o _ i [ 2 0 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 4   :   b e g i n  
                         p r i o _ i [ 2 1 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 8   :   b e g i n  
                         p r i o _ i [ 2 2 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 c   :   b e g i n  
                         p r i o _ i [ 2 3 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 0   :   b e g i n  
                         p r i o _ i [ 2 4 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 4   :   b e g i n  
                         p r i o _ i [ 2 5 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 8   :   b e g i n  
                         p r i o _ i [ 2 6 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 c   :   b e g i n  
                         p r i o _ i [ 2 7 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 0   :   b e g i n  
                         p r i o _ i [ 2 8 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 4   :   b e g i n  
                         p r i o _ i [ 2 9 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 2 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 8   :   b e g i n  
                         p r i o _ i [ 3 0 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         p r i o _ w e _ o [ 3 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 0 0   :   b e g i n  
                         i e _ i [ 0 ] [ 3 0 : 0 ]   =   r e q _ i . w d a t a [ 3 0 : 0 ] ;  
                         i e _ w e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 8 0   :   b e g i n  
                         i e _ i [ 1 ] [ 3 0 : 0 ]   =   r e q _ i . w d a t a [ 3 0 : 0 ] ;  
                         i e _ w e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   t h r e s h o l d  
                     3 2 ' h c 2 0 0 0 0 0   :   b e g i n  
                         t h r e s h o l d _ i [ 0 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         t h r e s h o l d _ w e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   t h r e s h o l d  
                     3 2 ' h c 2 0 1 0 0 0   :   b e g i n  
                         t h r e s h o l d _ i [ 1 ] [ 2 : 0 ]   =   r e q _ i . w d a t a [ 2 : 0 ] ;  
                         t h r e s h o l d _ w e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   c c  
                     3 2 ' h c 2 0 0 0 0 4   :   b e g i n  
                         c c _ i [ 0 ] [ 4 : 0 ]   =   r e q _ i . w d a t a [ 4 : 0 ] ;  
                         c c _ w e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   w r i t e   l o g i c   f o r   c c  
                     3 2 ' h c 2 0 1 0 0 4   :   b e g i n  
                         c c _ i [ 1 ] [ 4 : 0 ]   =   r e q _ i . w d a t a [ 4 : 0 ] ;  
                         c c _ w e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     d e f a u l t :   b e g i n    
                         r e s p _ o . e r r o r   =   1 ' b 1 ;  
                     e n d  
                 e n d c a s e  
             e n d   e l s e   b e g i n  
                 u n i q u e   c a s e ( r e q _ i . a d d r )  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 4   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 1 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 8   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 2 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 0 c   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 3 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 4 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 4   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 5 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 8   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 6 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 1 c   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 7 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 8 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 4   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 9 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 8   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 1 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 2 c   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 1 1 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 1 2 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 4   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 1 3 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 8   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 1 4 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 3 c   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 1 5 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 1 6 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 4   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 1 7 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 8   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 1 8 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 4 c   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 1 9 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 1 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 2 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 4   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 2 1 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 8   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 2 2 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 2 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 5 c   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 2 3 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 3 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 2 4 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 4 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 4   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 2 5 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 5 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 8   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 2 6 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 6 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 6 c   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 2 7 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 7 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 2 8 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 8 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 4   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 2 9 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 2 9 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   p r i o  
                     3 2 ' h c 0 0 0 0 7 8   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   p r i o _ o [ 3 0 ] [ 2 : 0 ] ;  
                         p r i o _ r e _ o [ 3 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i p  
                     3 2 ' h c 0 0 1 0 0 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 3 0 : 0 ]   =   i p _ o [ 3 0 : 0 ] ;  
                         i p _ r e _ o   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 0 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 3 0 : 0 ]   =   i e _ o [ 0 ] [ 3 0 : 0 ] ;  
                         i e _ r e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   i e  
                     3 2 ' h c 0 0 2 0 8 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 3 0 : 0 ]   =   i e _ o [ 1 ] [ 3 0 : 0 ] ;  
                         i e _ r e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   t h r e s h o l d  
                     3 2 ' h c 2 0 0 0 0 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   t h r e s h o l d _ o [ 0 ] [ 2 : 0 ] ;  
                         t h r e s h o l d _ r e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   t h r e s h o l d  
                     3 2 ' h c 2 0 1 0 0 0   :   b e g i n  
                         r e s p _ o . r d a t a [ 2 : 0 ]   =   t h r e s h o l d _ o [ 1 ] [ 2 : 0 ] ;  
                         t h r e s h o l d _ r e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   c c  
                     3 2 ' h c 2 0 0 0 0 4   :   b e g i n  
                         r e s p _ o . r d a t a [ 4 : 0 ]   =   c c _ o [ 0 ] [ 4 : 0 ] ;  
                         c c _ r e _ o [ 0 ]   =   1 ' b 1 ;  
                     e n d  
                     / /   r e a d   l o g i c   f o r   c c  
                     3 2 ' h c 2 0 1 0 0 4   :   b e g i n  
                         r e s p _ o . r d a t a [ 4 : 0 ]   =   c c _ o [ 1 ] [ 4 : 0 ] ;  
                         c c _ r e _ o [ 1 ]   =   1 ' b 1 ;  
                     e n d  
                     d e f a u l t :   b e g i n    
                         r e s p _ o . e r r o r   =   1 ' b 1 ;  
                     e n d  
                 e n d c a s e  
             e n d  
         e n d  
     e n d   :   e n d _ g e n _ r e g _ m u x _ p l i c _ r e g s  
 e n d m o d u l e  
  
 